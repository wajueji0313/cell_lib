module test_new (

);

endmodule
