module axis2axi (


);



endmodule 
