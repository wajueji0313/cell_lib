module test (

);


endmodule
