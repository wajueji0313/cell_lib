module test (

);
dsafasdgasgasgasgsagsa`1

endmodule
