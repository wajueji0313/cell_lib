module mem_ctrl(

):


endmodule
