module test_2 (



);


endmodule
